package metrics_pkg;

  import uvm_pkg::*;
 `include "uvm_macros.svh"

 `include "metric.sv"
 `include "metric_analyzer.sv"

endpackage: metrics_pkg
